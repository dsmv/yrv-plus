package tb_0_fabric_pkg;


class tb_0_fabric;

endclass
  
endpackage